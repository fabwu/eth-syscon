`timescale 1ns / 1ps // ETRM instruction memory 5.10.19
`default_nettype none

module IM #(parameter Inst=0, IAW=8, Size=256) (input wclk, rclk, wr, rd, input [IAW-1:0] wadr, radr,
      input wire [15:0] wdata, output wire [15:0] rdata);

wire [15:0] rdat [0:IAW-8];
if (IAW > 8) begin
	wire [IAW-9:0] bradr, bwadr;
	reg [IAW-9:0] bradrr;
	assign bwadr = wadr[IAW-1:8];
	assign bradr = radr[IAW-1:8];
	assign rdata = rdat[bradrr];
end
else
begin
	wire bradr;
	wire bwadr;
	reg bradrr;
	assign bradr = 0;
	assign bwadr = 0;
	assign rdata = rdat[0];
end


always @ (posedge rclk) begin
	if (rd)	
		bradrr <= bradr;
end

genvar i;
generate for (i = 0; i < Size / 256; i = i + 1) begin
SB_RAM40_4K #(.READ_MODE(0), .WRITE_MODE(0),
  .INIT_0(256'hFEEDC0DE0000000000000000000000000000000000000000FFFFD200C20F103F + (Inst << 192) + (i << 128)),
  .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
  .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000))
  bram(.WCLK(wclk), .RCLK(rclk), .WE(wr & (bwadr == i)), .RE(rd),
    .WCLKE(1'b1), .RCLKE(1'b1), .MASK(16'b0),
    .WADDR({3'b0, wadr[7:0]}), .RADDR({3'b0, radr[7:0]}), .WDATA(wdata), .RDATA(rdat[i]));
end endgenerate
endmodule

