`ifndef UtilityMacros_vh
`define UtilityMacros_vh

`define MAX(p,q) ((p)>(q)) ? (p) : (q)
`define MIN(p,q) ((p)<(q)) ? (p) : (q)

`endif